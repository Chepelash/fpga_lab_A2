module serializer_tb;




endmodule
